`pragma once

