import com_pkg::*;
`include "common/com_if.svh"

module rename(
    input clk,
    input rst,
    input clk_en,

    input flush_t flush,
    input stall,

    id3_rn_if.rename
);
    
endmodule
