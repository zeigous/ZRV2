import com_pkg::*;
`include "common/com_if.svh"

