module testbench (
    input clk,
    input clkEn,
    input rst
);
    
endmodule : testbench
